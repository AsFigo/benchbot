-- DUT file: ../examples/af_ud_counter/dut_src/af_up_dn_counter.vhdl
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;
use std.textio.all;
-- Adding OSVVM support below 
library osvvm;
context osvvm.OsvvmContext;

entity tb_af_up_dn_counter is

end entity tb_af_up_dn_counter;
