-- Generated using Python Parser for VHDL

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.numeric_std.all;
use std.textio.all;
-- User enabled --osvvm option 
-- Adding OSVVM support below 
library osvvm;
context osvvm.OsvvmContext;

entity tb_af_up_dn_counter is

end entity tb_af_up_dn_counter;
